entity full_adder is
  port (
    i_bit1  : in bit;
    i_bit2  : in bit;
    i_carry : in bit;
    --
    o_sum   : out bit;
    o_carry : out bit
  );
end full_adder;


architecture rtl of full_adder is

begin

end rtl;