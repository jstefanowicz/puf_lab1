entity adder4bit is
  port (
    i_in1     : in bit_vector(3 downto 0);
    i_in2     : in bit_vector(3 downto 0);
    --
    o_sum   : out bit_vector (3 downto 0);
    o_carry : out bit
  );
end adder4bit;


architecture rtl of adder4bit is


begin
  

  
end rtl;